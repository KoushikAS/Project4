module decoder5_32(i, o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31);
	input[4:0] i;
	output o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
	o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31;
	
	wire[4:0] n ;
	
	not n0(n[0],i[0]);
	not n1(n[1],i[1]);
	not n2(n[2],i[2]);
	not n3(n[3],i[3]);
	not n4(n[4],i[4]);
	
	
	and(o0, n[0],n[1], n[2], n[3], n[4]);
	and(o1, i[0],n[1], n[2], n[3], n[4]);
	and(o2, n[0],i[1], n[2], n[3], n[4]);
	and(o3, i[0],i[1], n[2], n[3], n[4]);
	and(o4, n[0],n[1], i[2], n[3], n[4]);
	and(o5, i[0],n[1], i[2], n[3], n[4]);
	and(o6, n[0],i[1], i[2], n[3], n[4]);
	and(o7, i[0],i[1], i[2], n[3], n[4]);
	and(o8, n[0],n[1], n[2], i[3], n[4]);
	and(o9, i[0],n[1], n[2], i[3], n[4]);
	and(o10, n[0],i[1], n[2], i[3], n[4]);
	and(o11, i[0],i[1], n[2], i[3], n[4]);
	and(o12, n[0],n[1], i[2], i[3], n[4]);
	and(o13, i[0],n[1], i[2], i[3], n[4]);
	and(o14, n[0],i[1], i[2], i[3], n[4]);
	and(o15, i[0],i[1], i[2], i[3], n[4]);
	and(o16, n[0],n[1], n[2], n[3], i[4]);
	and(o17, i[0],n[1], n[2], n[3], i[4]);
	and(o18, n[0],i[1], n[2], n[3], i[4]);
	and(o19, i[0],i[1], n[2], n[3], i[4]);
	and(o20, n[0],n[1], i[2], n[3], i[4]);
	and(o21, i[0],n[1], i[2], n[3], i[4]);
	and(o22, n[0],i[1], i[2], n[3], i[4]);
	and(o23, i[0],i[1], i[2], n[3], i[4]);
	and(o24, n[0],n[1], n[2], i[3], i[4]);
	and(o25, i[0],n[1], n[2], i[3], i[4]);
	and(o26, n[0],i[1], n[2], i[3], i[4]);
	and(o27, i[0],i[1], n[2], i[3], i[4]);
	and(o28, n[0],n[1], i[2], i[3], i[4]);
	and(o29, i[0],n[1], i[2], i[3], i[4]);
	and(o30, n[0],i[1], i[2], i[3], i[4]);
	and(o31, i[0],i[1], i[2], i[3], i[4]);
	
endmodule 